library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all ; 
use ieee.numeric_std.ALL;

entity breakout is
  port (    
    clk27M, reset_button      : in  std_logic;
	 SW								: in std_logic_vector(9 downto 0);
	 HEX0							   : out std_logic_vector(6 downto 0);
	 HEX1                      : out std_logic_vector(6 downto 0);
	 HEX2                      : out std_logic_vector(6 downto 0);
	 HEX3                      : out std_logic_vector(6 downto 0);
	 KEY                       : in std_logic_vector(3 downto 0);
	 LEDR                      : out std_logic_vector(9 downto 0);
	 LEDG                      : out std_logic_vector(7 downto 0);
    red, green, blue          : out std_logic_vector(3 downto 0);
    hsync, vsync              : out std_logic);
end breakout;

architecture comportamento of breakout is
 
  component ball
	port (clk27M		 : in std_logic;
		rstn 		    	 : in std_logic;
		paddle_size     : in integer range 0 to 10;
		paddle_X		    : in integer range 0 to 128;
		paddle_Y	   	 : in integer range 0 to 95;
		ball_X    		 : buffer integer range 0 to 128;
		ball_Y	   	 : buffer integer range 0 to 95;
		colision		    : in std_logic;
		trapaca			 : in std_logic;
		speed_control   : in std_logic);
  
  end component;
  
	component brick
		port (clk27M	 : in std_logic;
			rstn 			 : in std_logic;
			ball_X		 : in integer range 0 to 128;
			ball_Y		 : in integer range 0 to 95;
			colision 	 : out std_logic;
			condition    : buffer std_logic_vector (128 downto 0);
			condition2   : buffer std_logic_vector (128 downto 0);
			condition3   : buffer std_logic_vector (128 downto 0));
	end component;
	
	component contador_pontos
	PORT ( 	Clock 								: in std_logic;
				Enable 								: in std_logic;
				n_pontos 						   : in integer range 0 to 128;
				Clear									: IN STD_LOGIC;
				BCD3, BCD2, BCD1, BCD0	 		: BUFFER  STD_LOGIC_VECTOR(3 DOWNTO 0)
				);
	end component;
	
	component display7seg
	port (Inp : in std_logic_vector(3 downto 0);
			Xis : out std_logic_vector(6 downto 0)
	);		  

	end component;

	component controle_pontos
		port (clk27M				 : in std_logic;
		rstn 	    					 : in std_logic;
		colision  	           	 : in std_logic;
		jogo_start 	         	 : in std_logic;
		ball_Y			  	 		 : in integer range 0 to 95;
		LEDR 							 : out std_logic_vector(9 downto 0); 
		reset_ball 				    : out std_logic; 
		reset_brick					 : out std_logic;
		speed_control 				 : out std_logic;
		game_over_control        : out std_logic;
		win_game_control 			 : out std_logic;
		brick_condition          : in std_logic_vector (128 downto 0);
		brick_condition2 			 : in std_logic_vector(128 downto 0);
		brick_condition3 			 : in std_logic_vector(128 downto 0);
		n_pontos 					 : out integer range 0 to 128;
		trapaca   					 : in std_logic
		);
	end component;

  signal rstn : std_logic;  -- reset active low

  -- Interface com a memoria de video
  signal we : std_logic;                        -- write enable ('1' p/ escrita)
  signal addr : integer range 0 to 12287;       -- endereco mem. vga
  signal pixel : std_logic_vector(2 downto 0);  -- valor de cor do pixel
  signal pixel_bit : std_logic;                 -- um bit do vetor acima
  
  -- Sinais dos contadores de linhas e colunas utilizados para percorrer
  -- as posicoes da memoria de video (pixels) no momento de construir um quadro.
  
  signal line : integer range 0 to 95;  -- linha atual
  signal col : integer range 0 to 127;  -- coluna atual

  signal col_rstn : std_logic;          -- reset do contador de colunas
  signal col_enable : std_logic;        -- enable do contador de colunas

  signal line_rstn : std_logic;          -- reset do contador de linhas
  signal line_enable : std_logic;        -- enable do contador de linhas

  signal fim_escrita : std_logic;       -- '1' quando um quadro terminou de ser escrito 


  --sinais para a posicao da raquete
  signal pos_x : integer range 0 to 127;
  signal pos_y : integer range 0 to 95;
  
  signal atualiza_pos_x : std_logic;    -- se '1' = bola muda sua pos. no eixo x
  
	--sinais que armazenam a posicao da nossa bolinha
	signal ball_X : integer range 0 to 127;
	signal ball_Y : integer range 0 to 95;

	--sinais para controlar quais tijolos ja foram quebrados
	signal brick_condition : std_logic_vector (128 downto 0);
	signal brick_condition2 : std_logic_vector (128 downto 0);
	signal brick_condition3 : std_logic_vector (128 downto 0);
	
	--sinal para controlar nossos pontos
	signal n_pontos :  integer range 0 to 128;
	
  -- Tipos e sinais da maquina de estados de controle
  type estado_t is (show_splash, inicio, constroi_quadro, move_bola);
  signal estado: estado_t := show_splash;
  signal proximo_estado: estado_t := show_splash;

  --sinais para o um contador para controlarmos a velocidade
  --de atualizacao da posicao do paddle
  signal contador : integer range 0 to 270000 - 1;  -- contador
  signal timer : std_logic;        -- vale '1' quando o contador chegar ao fim
  signal timer_rstn, timer_enable : std_logic;
  
  
  --constante para o tamanho da raquete
  constant paddle_size : integer := 10;
  
  --sinal que indica colisao da bola com um tijolo
  signal colision : std_logic;
  
  --sinal para resetarmos apenas a posicao da bola
  signal reset_ball : std_logic;
  
  --sinal para resetarmos apenas os tijolos (reconstruir)
  signal reset_brick : std_logic;
  
  --sinais para fim de jogo e comeco de jogo
  signal game_over_control  : std_logic;
  signal win_game_control   : std_logic;
  
  --flag para alternar entre as duas velocidade da bola
  signal speed_control : std_logic;

  --sinais para os contadores
  signal BCD0 : std_logic_vector (3 downto 0);
  signal BCD1 : std_logic_vector (3 downto 0);
  signal BCD2 : std_logic_vector (3 downto 0);
  signal BCD3 : std_logic_vector (3 downto 0);
  
  --sprites
  signal game_over_sprite : std_logic_vector (12192 downto 0);
  signal win_game_sprite  : std_logic_vector (12192 downto 0);
  
begin  -- comportamento

  --instancia nossa bolinha
	ball_inst : ball port map (clk27M, reset_ball, paddle_size, pos_x, pos_y, ball_X, ball_Y, colision, SW(8), speed_control);
  
	
	--instancia o gerenciador dos tijolos
	brick_gen : brick port map (clk27M, reset_brick, ball_X, ball_Y, colision,brick_condition (128 downto 0), brick_condition2(128 downto 0), brick_condition3(128 downto 0));  
  
   --instancia o controlador de pontos e fase
	controle_inst : controle_pontos port map (clk27M, rstn, colision, KEY(1), ball_Y ,LEDR(9 downto 0), reset_ball, reset_brick, speed_control, game_over_control, win_game_control ,brick_condition(128 downto 0), brick_condition2(128 downto 0), brick_condition3(128 downto 0), n_pontos, SW(9));
  
	--instancia o contador de pontos
	cont_pont_inst : contador_pontos port map (clk27M, colision , n_pontos, rstn, BCD3(3 downto 0), BCD2(3 downto 0), BCD1(3 downto 0),BCD0(3 downto 0));
	
	--instancia os display7seg
	display1_inst : display7seg port map (BCD0(3 downto 0), HEX0(6 downto 0));
	display2_inst : display7seg port map (BCD1(3 downto 0), HEX1(6 downto 0));
	display3_inst : display7seg port map (BCD2(3 downto 0), HEX2(6 downto 0));
	display4_inst : display7seg port map (BCD3(3 downto 0), HEX3(6 downto 0));
	
  -- Instancia do controlador de video: 128 colunas por 96 linhas
  -- (aspect ratio 4:3). Os sinais que iremos utilizar para comunicar
  -- com a memoria de video (para alterar o brilho dos pixels) sao
  -- write_clk (nosso clock), write_enable ('1' quando queremos escrever
  -- o valor de um pixel), write_addr (endereco do pixel a escrever)
  -- e data_in (valor do brilho do pixel RGB, 1 bit pra cada componente de cor)
	vga_controller: entity work.vgacon port map (
		clk27M       => clk27M,
		rstn         => '1',
		red          => red,
		green        => green,
		blue         => blue,
		hsync        => hsync,
		vsync        => vsync,
		write_clk    => clk27M,
		write_enable => we,
		write_addr   => addr,
		data_in      => pixel);
	
  --percorre todas as linhas e colunas desenhando o quadro do jogo
  conta_coluna: process (clk27M, col_rstn)
  begin 
    if col_rstn = '0' then                  
      col <= 0;
    elsif clk27M'event and clk27M = '1' then
      if col_enable = '1' then
        if col = 127 then   
          col <= 0;
        else
          col <= col + 1;  
        end if;
      end if;
    end if;
  end process conta_coluna;

  conta_linha: process (clk27M, line_rstn)
  begin  
    if line_rstn = '0' then                 
      line <= 0;
    elsif clk27M'event and clk27M = '1' then  
      --passa de linha depois de contar todas as colunas
      if line_enable = '1' and col = 127 then
        if line = 95 then   -- conta de 0 a 95 (96 linhas)
          line <= 0;
        else
          line <= line + 1;  
        end if;        
      end if;
    end if;
  end process conta_linha;

   --indica que o quadro ja foi construido
   fim_escrita <= '1' when (line = 95) and (col = 127)  else '0';   
   
	--esse processo autaliza a posicao da raquete
	p_atualiza_pos_x: process (clk27M, rstn)
	--contador para termos 60Hz de taxa de atualizacao
	variable contador : integer range 0 to 450000;
	
	begin 
    if rstn = '0' then                  
      pos_x <= 64;		 --posicao da raquete					 
		pos_y <= 80;							 
		contador := 0;
		
    elsif clk27M'event and clk27M = '1' then
      contador := contador + 1;
		
		--contador para atualizarmos a posicao em velocidade adequada
		if contador >= 449999 then
		  contador := 0;
			
		  --muda a posicao da raquete de acordo com os inputs
        if KEY(2) = '0' then         
			 --nao deixa a raquete ultrapassar as bordas
          if (pos_x+paddle_size) = 127 then
            pos_x <= pos_x;  
				
          else
				--move a raquete
            pos_x <= pos_x + 1;
		   end if;        
			
			elsif KEY(3) = '0' then
				--nao deixa a raquete ultrapassar as bordas
				if (pos_x-paddle_size) = 0 then
					pos_x <= pos_x;
          
				else
					--move a raquete
					pos_x <= pos_x - 1;
				end if;
			end if;
		end if;
	end if;
  end process p_atualiza_pos_x;


	--sprites de game over e de win game
	game_over_sprite <= "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111110000000000000000111000000000000001100000000000011100000001111111111111111111111100000000000000000000000000000000001100000000000000000000000000110110000000000000111000000000011110000000111111111111111111111110000000000000000000000000000000000110000000000000000000000000110001100000000000011011000000011011000000011100000000000000000000000000000000000000000000000000000011000000000000000000000000110000011000000000001100110000011001100000001110000000000000000000000000000000000000000000000000000001100000000000000000000001110000000110000000000110001100011000110000000111000000000000000000000000000000000000000000000000000000110000111111111100000001110000000001100000000011000011011000011000000011111111111111111111111000000000000000000000000000000000011000011111111110000000110000000000011000000001100000111000001100000001111111111111111111111100000000000000000000000000000000001100000000000011000000111111111111111110000000110000001000000110000000111000000000000000000000000000000000000000000000000000000110000000000001100000111111111111111111100000011000000000000011000000011100000000000000000000000000000000000000000000000000000011000000000000110000110000000000000000011000001100000000000001100000001110000000000000000000000000000000000000000000000000000001100000000000011000110000000000000000000110000110000000000000110000000111111111111111111111110000000000000000000000000000000000111111111111111100110000000000000000000001100011000000000000011000000011111111111111111111111000000000000000000000000000000000011111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111110010000000000000000000000000100000111111111111111111111000000000111111111111000000000000000000000000000000000000010000000000001000100000000000000000000000100000010000000000000000000000000000010000000000010000000000000000000000000000000000001000000000000100001000000000000000000000100000001000000000000000000000000000001000000000000100000000000000000000000000000000000100000000000010000010000000000000000000100000000100000000000000000000000000000100000000000001000000000000000000000000000000000010000000000001000000100000000000000000100000000010000000000000000000000000000010000000000000100000000000000000000000000000000001000000000000100000001000000000000000100000000001000000000000000000000000000001000000000000010000000000000000000000000000000000100000000000010000000010000000000000100000000000111111111111111111111000000000111111111111110000000000000000000000000000000000010000000000001000000000100000000000100000000000010000000000000000000000000000011000000000000000000000000000000000000000000000001000000000000100000000001000000000100000000000001000000000000000000000000000001010000000000000000000000000000000000000000000000100000000000010000000000010000000100000000000000100000000000000000000000000000100100000000000000000000000000000000000000000000010000000000001000000000000100000100000000000000010000000000000000000000000000010001000000000000000000000000000000000000000000001000000000000100000000000001000100000000000000001000000000000000000000000000001000011000000000000000000000000000000000000000000100000000000010000000000000010100000000000000000100000000000000000000000000000100000011000000000000000000000000000000000000000011111111111111000000000000000100000000000000000011111111111111111111100000000010000000011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	win_game_sprite  <= "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100000000000000000011000000000111111111111111111111111110000000001100000000000000110000000000000000000000000000000000000000000011000000000000000011000000000011111111111111111111111111000000000110000000000000011000000000000000000000000000000000000000000000011000000000000011000000000001110000000000000000000011100000000011000000000000001100000000000000000000000000000000000000000000000110000000000011000000000000111000000000000000000001110000000001100000000000000110000000000000000000000000000000000000000000000001100000000011000000000000011100000000000000000000111000000000110000000000000011000000000000000000000000000000000000000000000000011100000011000000000000001110000000000000000000011100000000011000000000000001100000000000000000000000000000000000000000000000000011000011000000000000000111000000000000000000001110000000001100000000000000110000000000000000000000000000000000000000000000000000110011000000000000000011100000000000000000000111000000000110000000000000011000000000000000000000000000000000000000000000000000000111000000000000000001110000000000000000000011100000000011000000000000001100000000000000000000000000000000000000000000000000000011100000000000000000111000000000000000000001110000000001100000000000000110000000000000000000000000000000000000000000000000000001110000000000000000011100000000000000000000111000000000110000000000000011000000000000000000000000000000000000000000000000000000111000000000000000001110000000000000000000011100000000011000000000000001100000000000000000000000000000000000000000000000000000011100000000000000000111000000000000000000001110000000001100000000000000110000000000000000000000000000000000000000000000000000001110000000000000000011100000000000000000000111000000000110000000000000110000000000000000000000000000000000000000000000000000000111000000000000000001110000000000000000000011100000000001100000000000110000000000000000000000000000000000000000000000000000000011100000000000000000111111111111111111111111110000000000011111111111110000000000000000000000000000000000000000000000000000000001110000000000000000011111111111111111111111111000000000000111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110000000000001110000000000110000000001111111111111111111111111000000111111000000000000111000000000000000000000000000000000000001110000000000111000000000110000000000111111111111111111111111100000011111110000000000011100000000000000000000000000000000000000011100000000011100000000011000000000011000000000000000000000110000001110011110000000001110000000000000000000000000000000000000000110000000001110000000011100000000001100000000000000000000011000000111000011100000000111000000000000000000000000000000000000000001100000000111000000001100000000000110000000000000000000001100000011100000111000000011100000000000000000000000000000000000000000110000000011100000000110000000000011000000000000000000000110000001110000001110000001110000000000000000000000000000000000000000011100000001110000000011000000000001100000000000000000000011000000111000000011100000111000000000000000000000000000000000000000000110000000111000000011100000000000110000000000000000000001100000011100000000111000011100000000000000000000000000000000000000000011000000011100000001110000000000011000000000000000000000110000001110000000001110001110000000000000000000000000000000000000000001110000001110000001110000000000001100000000000000000000011000000111000000000011100111000000000000000000000000000000000000000000111000000111000001110000000000000110000000000000000000001100000011100000000000110110000000000000000000000000000000000000000000000111111111111111100000000000000011111111111111111111111110000001110000000000001111000000000000000000000000000000000000000000000011111111111111110000000000000001111111111111111111111111000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111110000000000000000000000000000000000001111111111000000000000000000000000000000000000000000000000000000000000000000000011000000011000000000000000000000000000000000000110000001100000000000000000000000000000000000000000000000000000000000000000000011100000011110000000000000000000000000000000000111000000111000000000000000000000000000000000000000000000000000000000000000000000110000000110000000000000000000000000000000000001100000011000000000000000000000000000000000000000000000000000000000000000000000011000000011000000000000000000000000000000000000111111111100000000000000000000000000000000000000000000000000000000000000000000001111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000010000000000010000000010000000100000001000000000110000000000000000000000000000000000000000000000000000000000000000000000000000001110000000001000000001000000010000000100000000110000000000000000000000000000000000000000000000000000000000000000000000000000000001110000000100000000100000001000000010000000110000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110000000100000010000001000000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110000001000000100000100000000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110000100000010000010000001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
  
	--desenha os pixels na tela
	pixel_process:	process (clk27M, rstn)
	begin
		--desenha a tela de game over, se for o caso
		if(game_over_control = '1') then
			if (game_over_sprite((96 - line)*127 + (127 - col)) = '1') then
				pixel <= "101";
				
			else
				pixel <= "000";
			end if;
		
		--desenha a tela de win game, se for o caso
		elsif (win_game_control = '1') then
			if (win_game_sprite((96 - line)*127 + (127 - col)) = '1') then
				pixel <= "101";
				
			else
				pixel <= "000";
			end if;
		
		--desenha a raquete
		elsif((col <= pos_x + paddle_size) and (col >= pos_x - paddle_size) and (line = pos_y)) then
			pixel <= "111";
		
		--desenha a bolinha
		elsif	( (col = ball_X) and (line = ball_Y) ) then
		pixel <= "111";
		
		--desenha a primeira barra de tijolos
		elsif (line = 5 OR line = 6 OR line = 7 or line = 8 OR line = 9 OR line = 10 OR line = 11 or line = 12 )		then
			--percorre todas as colunas
			for I in 0 to 127 loop 
				if (brick_condition(I) = '1' and col = I) then
					pixel <= "011";
					
				elsif(brick_condition(I) = '0' and col = I) then
					pixel <= "000";
				end if;
			end loop;
			
		--desenha a segunda barra de tijolos
		elsif (line = 13 OR line = 14 OR line = 15 OR line = 16 OR line = 17 OR line = 18 OR line = 19 OR line = 20) then
			--percorre todas as colunas
			for I in 0 to 127 loop 
				if (brick_condition2(I) = '1' and col = I) then
					pixel <= "001";
					
				elsif(brick_condition2(I) = '0' and col = I) then
					pixel <= "000";
				end if;
			end loop;
			
		--desenha a terceira barra de tijolos
		elsif (line = 21 OR line = 22 OR line = 23 OR line = 24 OR line = 25 OR line = 26 OR line = 27 OR line = 28) then
			--percorre todas as colunas
			for I in 0 to 127 loop 
				if (brick_condition3(I) = '1' and col = I) then
					pixel <= "110";
					
				elsif(brick_condition3(I) = '0' and col = I) then
					pixel <= "000";
				end if;
			end loop;
			
		--deixa preto os outros pixels
		else
			pixel <= "000";
			
		end if;
		
	end process pixel_process;
	 
  --endereco da memoria
  addr  <= col + (128 * line);

  --processo para a maquina de estado de controle
  logica_mealy: process (estado, fim_escrita, timer)
  begin 
    case estado is
      when inicio         => if timer = '1' then              
                               proximo_estado <= constroi_quadro;
                             else
                               proximo_estado <= inicio;
                             end if;
                             atualiza_pos_x <= '0';
                             line_rstn      <= '0';  -- reset � active low!
                             line_enable    <= '0';
                             col_rstn       <= '0';  -- reset � active low!
                             col_enable     <= '0';
                             we             <= '0';
                             timer_rstn     <= '1';  -- reset � active low!
                             timer_enable   <= '1';

      when constroi_quadro=> if fim_escrita = '1' then
                               proximo_estado <= move_bola;
                             else
                               proximo_estado <= constroi_quadro;
                             end if;
                             atualiza_pos_x <= '0';
                             line_rstn      <= '1';
                             line_enable    <= '1';
                             col_rstn       <= '1';
                             col_enable     <= '1';
                             we             <= '1';
                             timer_rstn     <= '0'; 
                             timer_enable   <= '0';

      when move_bola      => proximo_estado <= inicio;
                             atualiza_pos_x <= '1';
                             line_rstn      <= '1';
                             line_enable    <= '0';
                             col_rstn       <= '1';
                             col_enable     <= '0';
                             we             <= '0';
                             timer_rstn     <= '0'; 
                             timer_enable   <= '0';

      when others         => proximo_estado <= inicio;
                             atualiza_pos_x <= '0';
                             line_rstn      <= '1';
                             line_enable    <= '0';
                             col_rstn       <= '1';
                             col_enable     <= '0';
                             we             <= '0';
                             timer_rstn     <= '1'; 
                             timer_enable   <= '0';
      
    end case;
  end process logica_mealy;
  
  --muda o estado da maquina de estado
  seq_fsm: process (clk27M, rstn)
  begin 
    if rstn = '0' then
      estado <= inicio;
    elsif clk27M'event and clk27M = '1' then 
      estado <= proximo_estado;
    end if;
  end process seq_fsm;

 
  --contador para termos os 60Hz a partir do clck da placa
  p_contador: process (clk27M, timer_rstn)
  begin
    if timer_rstn = '0' then     
      contador <= 0;
    elsif clk27M'event and clk27M = '1' then  
      if timer_enable = '1' then       
        if contador = 270000 - 1 then
          contador <= 0;
        else
          contador <=  contador + 1;        
        end if;
      end if;
    end if;
  end process p_contador;

 
  --indica que nosso contador terminou de contar
  p_timer: process (contador)
  begin
    if contador = 270000 - 1 then
      timer <= '1';
    else
      timer <= '0';
    end if;
  end process p_timer;

  -----------------------------------------------------------------------------
  -- Processos que sincronizam sinais assincronos, de preferencia com mais
  -- de 1 flipflop, para evitar metaestabilidade.
  -----------------------------------------------------------------------------
  
  -- purpose: Aqui sincronizamos nosso sinal de reset vindo do botao da DE1
  -- type   : sequential
  -- inputs : clk27M
  -- outputs: rstn
  build_rstn: process (clk27M)
		variable temp : std_logic;          -- flipflop intermediario
  begin  
		if clk27M'event and clk27M = '1' then 
			rstn <= temp;
			temp := reset_button;      
    end if;
  end process build_rstn;
  
end comportamento;
